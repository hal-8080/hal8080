LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY main_memory IS
	PORT(
		
	);
END ENTITY main_memory;
ARCHITECTURE bhv OF main_memory IS

BEGIN

END;