--             HAL8080 Processor           --
-- Dennis, Kasper, Tjeerd, Nick, Oussama 2020
--                control
-- The processor control.

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY control IS
    PORT(
        clk : IN std_logic -- Main (50Mhz) clock.
    );
END ENTITY control;

ARCHITECTURE bhv OF control IS
BEGIN

END bhv;