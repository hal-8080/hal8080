--             HAL8080 Processor           --
-- Dennis, Kasper, Tjeerd, Nick, Oussama 2020
--                memory
-- This file describes the hardware for the main
-- memory.

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY memory IS
    PORT (
        clk : IN std_logic -- Main (50Mhz) clock.
    );
END ENTITY memory;

ARCHITECTURE bhv OF memory IS
BEGIN

END bhv;