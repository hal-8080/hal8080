--             HAL8080 Processor           --
-- Dennis, Kasper, Tjeerd, Nick, Oussama 2020
--                datapath
-- The processor datapath.

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY datapath IS
    PORT(
        clk : IN std_logic -- Main (50Mhz) clock.
    );
END ENTITY datapath;

ARCHITECTURE bhv OF datapath IS
BEGIN

END bhv;